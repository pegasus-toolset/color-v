module color

pub struct Color {
pub:
	r byte
	g byte
	b byte
	a byte = byte(255)
}

pub const (
	// Pink colors
	pink              = Color{r: 0xFF, g: 0xC0, b: 0xCB}
	light_pink        = Color{r: 0xFF, g: 0xB6, b: 0xC1}
	hot_pink          = Color{r: 0xFF, g: 0x69, b: 0xB4}
	deep_pink         = Color{r: 0xFF, g: 0x14, b: 0x93}
	pale_violet_red   = Color{r: 0xDB, g: 0x70, b: 0x93}
	medium_violet_red = Color{r: 0xC7, g: 0x15, b: 0x85}

	// Red colors
	light_salmon = Color{r: 0xFF, g: 0xA0, b: 0x7A}
	salmon       = Color{r: 0xFA, g: 0x80, b: 0x72}
	dark_salmon  = Color{r: 0xE9, g: 0x96, b: 0x7A}
	light_coral  = Color{r: 0xF0, g: 0x80, b: 0x80}
	indian_red   = Color{r: 0xCD, g: 0x5C, b: 0x5C}
	crimson      = Color{r: 0xDC, g: 0x14, b: 0x3C}
	firebrick    = Color{r: 0xB2, g: 0x22, b: 0x22}
	dark_red     = Color{r: 0x8B, g: 0x00, b: 0x00}
	red          = Color{r: 0xFF, g: 0x00, b: 0x00}

	// Orange colors
	orange_red  = Color{r: 0xFF, g: 0x45, b: 0x00}
	tomato      = Color{r: 0xFF, g: 0x63, b: 0x47}
	coral       = Color{r: 0xFF, g: 0x7F, b: 0x50}
	dark_orange = Color{r: 0xFF, g: 0x8C, b: 0x00}
	orange      = Color{r: 0xFF, g: 0xA5, b: 0x00}

	// Yellow colors
	yellow                 = Color{r: 0xFF, g: 0xFF, b: 0x00}
	light_yellow           = Color{r: 0xFF, g: 0xFF, b: 0xE0}
	lemon_chiffon          = Color{r: 0xFF, g: 0xFA, b: 0xCD}
	light_goldenrod_yellow = Color{r: 0xFA, g: 0xFA, b: 0xD2}
	papaya_whip            = Color{r: 0xFF, g: 0xEF, b: 0xD5}
	moccasin               = Color{r: 0xFF, g: 0xE4, b: 0xB5}
	peach_puff             = Color{r: 0xFF, g: 0xDA, b: 0xB9}
	pale_goldenrod         = Color{r: 0xEE, g: 0xE8, b: 0xAA}
	khaki                  = Color{r: 0xF0, g: 0xE6, b: 0x8C}
	dark_khaki             = Color{r: 0xBD, g: 0xB7, b: 0x6B}
	gold                   = Color{r: 0xFF, g: 0xD7, b: 0x00}

	// Brown colors
	cornsilk        = Color{r: 0xFF, g: 0xF8, b: 0xDC}
	blanched_almond = Color{r: 0xFF, g: 0xEB, b: 0xCD}
	bisque          = Color{r: 0xFF, g: 0xE4, b: 0xC4}
	navajo_white    = Color{r: 0xFF, g: 0xDE, b: 0xAD}
	wheat           = Color{r: 0xF5, g: 0xDE, b: 0xB3}
	burlywood       = Color{r: 0xDE, g: 0xB8, b: 0x87}
	tan             = Color{r: 0xD2, g: 0xB4, b: 0x8C}
	rosy_brown      = Color{r: 0xBC, g: 0x8F, b: 0x8F}
	sandy_brown     = Color{r: 0xF4, g: 0xA4, b: 0x60}
	goldenrod       = Color{r: 0xDA, g: 0xA5, b: 0x20}
	dark_goldenrod  = Color{r: 0xB8, g: 0x86, b: 0x0B}
	peru            = Color{r: 0xCD, g: 0x85, b: 0x3F}
	chocolate       = Color{r: 0xD2, g: 0x69, b: 0x1E}
	saddle_brown    = Color{r: 0x8B, g: 0x45, b: 0x13}
	sienna          = Color{r: 0xA0, g: 0x52, b: 0x2D}
	brown           = Color{r: 0xA5, g: 0x2A, b: 0x2A}
	maroon          = Color{r: 0x80, g: 0x00, b: 0x00}

	// Green colors
	dark_olive_green    = Color{r: 0x55, g: 0x6B, b: 0x2F}
	olive               = Color{r: 0x80, g: 0x80, b: 0x00}
	olive_drab          = Color{r: 0x6B, g: 0x8E, b: 0x23}
	yellow_green        = Color{r: 0x9A, g: 0xCD, b: 0x32}
	lime_green          = Color{r: 0x32, g: 0xCD, b: 0x32}
	lime                = Color{r: 0x00, g: 0xFF, b: 0x00}
	lawn_green          = Color{r: 0x7C, g: 0xFC, b: 0x00}
	chartreuse          = Color{r: 0x7F, g: 0xFF, b: 0x00}
	green_yellow        = Color{r: 0xAD, g: 0xFF, b: 0x2F}
	spring_green        = Color{r: 0x00, g: 0xFF, b: 0x7F}
	medium_spring_green = Color{r: 0x00, g: 0xFA, b: 0x9A}
	light_green         = Color{r: 0x90, g: 0xEE, b: 0x90}
	pale_green          = Color{r: 0x98, g: 0xFB, b: 0x98}
	dark_sea_green      = Color{r: 0x8F, g: 0xBC, b: 0x8F}
	medium_aquamarine   = Color{r: 0x66, g: 0xCD, b: 0xAA}
	medium_sea_green    = Color{r: 0x3C, g: 0xB3, b: 0x71}
	sea_green           = Color{r: 0x2E, g: 0x8B, b: 0x57}
	forest_green        = Color{r: 0x22, g: 0x8B, b: 0x22}
	green               = Color{r: 0x00, g: 0x80, b: 0x00}
	dark_green          = Color{r: 0x00, g: 0x64, b: 0x00}

	// Cyan colors
	aqua             = Color{r: 0x00, g: 0xFF, b: 0xFF}
	cyan             = Color{r: 0x00, g: 0xFF, b: 0xFF}
	light_cyan       = Color{r: 0xE0, g: 0xFF, b: 0xFF}
	pale_turquoise   = Color{r: 0xAF, g: 0xEE, b: 0xEE}
	aquamarine       = Color{r: 0x7F, g: 0xFF, b: 0xD4}
	turquoise        = Color{r: 0x40, g: 0xE0, b: 0xD0}
	medium_turquoise = Color{r: 0x48, g: 0xD1, b: 0xCC}
	dark_turquoise   = Color{r: 0x00, g: 0xCE, b: 0xD1}
	light_sea_green  = Color{r: 0x20, g: 0xB2, b: 0xAA}
	cadet_blue       = Color{r: 0x5F, g: 0x9E, b: 0xA0}
	dark_cyan        = Color{r: 0x00, g: 0x8B, b: 0x8B}
	teal             = Color{r: 0x00, g: 0x80, b: 0x80}

	// Blue colors
	light_steel_blue = Color{r: 0xB0, g: 0xC4, b: 0xDE}
	powder_blue      = Color{r: 0xB0, g: 0xE0, b: 0xE6}
	light_blue       = Color{r: 0xAD, g: 0xD8, b: 0xE6}
	sky_blue         = Color{r: 0x87, g: 0xCE, b: 0xEB}
	light_sky_blue   = Color{r: 0x87, g: 0xCE, b: 0xFA}
	deep_sky_blue    = Color{r: 0x00, g: 0xBF, b: 0xFF}
	dodger_blue      = Color{r: 0x1E, g: 0x90, b: 0xFF}
	cornflower_blue  = Color{r: 0x64, g: 0x95, b: 0xED}
	steel_blue       = Color{r: 0x46, g: 0x82, b: 0xB4}
	royal_blue       = Color{r: 0x41, g: 0x69, b: 0xE1}
	blue             = Color{r: 0x00, g: 0x00, b: 0xFF}
	medium_blue      = Color{r: 0x00, g: 0x00, b: 0xCD}
	dark_blue        = Color{r: 0x00, g: 0x00, b: 0x8B}
	navy             = Color{r: 0x00, g: 0x00, b: 0x80}
	midnight_blue    = Color{r: 0x19, g: 0x19, b: 0x70}

	// Purple, violet, and magenta colors
	lavender          = Color{r: 0xE6, g: 0xE6, b: 0xFA}
	thistle           = Color{r: 0xD8, g: 0xBF, b: 0xD8}
	plum              = Color{r: 0xDD, g: 0xA0, b: 0xDD}
	violet            = Color{r: 0xEE, g: 0x82, b: 0xEE}
	orchid            = Color{r: 0xDA, g: 0x70, b: 0xD6}
	fuchsia           = Color{r: 0xFF, g: 0x00, b: 0xFF}
	magenta           = Color{r: 0xFF, g: 0x00, b: 0xFF}
	medium_orchid     = Color{r: 0xBA, g: 0x55, b: 0xD3}
	medium_purple     = Color{r: 0x93, g: 0x70, b: 0xDB}
	blue_violet       = Color{r: 0x8A, g: 0x2B, b: 0xE2}
	dark_violet       = Color{r: 0x94, g: 0x00, b: 0xD3}
	dark_orchid       = Color{r: 0x99, g: 0x32, b: 0xCC}
	dark_magenta      = Color{r: 0x8B, g: 0x00, b: 0x8B}
	purple            = Color{r: 0x80, g: 0x00, b: 0x80}
	indigo            = Color{r: 0x4B, g: 0x00, b: 0x82}
	dark_slate_blue   = Color{r: 0x48, g: 0x3D, b: 0x8B}
	slate_blue        = Color{r: 0x6A, g: 0x5A, b: 0xCD}
	medium_slate_blue = Color{r: 0x7B, g: 0x68, b: 0xEE}

	// White colors
	white          = Color{r: 0xFF, g: 0xFF, b: 0xFF}
	snow           = Color{r: 0xFF, g: 0xFA, b: 0xFA}
	honeydew       = Color{r: 0xF0, g: 0xFF, b: 0xF0}
	mint_cream     = Color{r: 0xF5, g: 0xFF, b: 0xFA}
	azure          = Color{r: 0xF0, g: 0xFF, b: 0xFF}
	alice_blue     = Color{r: 0xF0, g: 0xF8, b: 0xFF}
	ghost_white    = Color{r: 0xF8, g: 0xF8, b: 0xFF}
	white_smoke    = Color{r: 0xF5, g: 0xF5, b: 0xF5}
	seashell       = Color{r: 0xFF, g: 0xF5, b: 0xEE}
	beige          = Color{r: 0xF5, g: 0xF5, b: 0xDC}
	old_lace       = Color{r: 0xFD, g: 0xF5, b: 0xE6}
	floral_white   = Color{r: 0xFF, g: 0xFA, b: 0xF0}
	ivory          = Color{r: 0xFF, g: 0xFF, b: 0xF0}
	antique_white  = Color{r: 0xFA, g: 0xEB, b: 0xD7}
	linen          = Color{r: 0xFA, g: 0xF0, b: 0xE6}
	lavender_blush = Color{r: 0xFF, g: 0xF0, b: 0xF5}
	misty_rose     = Color{r: 0xFF, g: 0xE4, b: 0xE1}

	// Gray and black colors
	gainsboro        = Color{r: 0xDC, g: 0xDC, b: 0xDC}
	light_gray       = Color{r: 0xD3, g: 0xD3, b: 0xD3}
	silver           = Color{r: 0xC0, g: 0xC0, b: 0xC0}
	dark_gray        = Color{r: 0xA9, g: 0xA9, b: 0xA9}
	gray             = Color{r: 0x80, g: 0x80, b: 0x80}
	dim_gray         = Color{r: 0x69, g: 0x69, b: 0x69}
	light_slate_gray = Color{r: 0x77, g: 0x88, b: 0x99}
	slate_gray       = Color{r: 0x70, g: 0x80, b: 0x90}
	dark_slate_gray  = Color{r: 0x2F, g: 0x4F, b: 0x4F}
	black            = Color{r: 0x00, g: 0x00, b: 0x00}
)

// equals return true if te given color is exactly equal to this color.
pub fn (this Color) equals(c Color) bool {
	return this.r == c.r && this.g == c.g && this.b == c.b && this.a == c.a
}

